
 module credit_bitmap (

	input	logic	clk, 
	input	logic	resetN, 
	input logic	[10:0] offsetX,// offset from top left  position 
	input logic	[10:0] offsetY, 
	input	logic	InsideRectangle, //input that the pixel is within a bracket 

	output	logic	drawingRequest, //output that the pixel should be dispalyed 
	output	logic	[11:0] RGBout,  //rgb value from the bitmap 
	output	logic	[3:0] HitEdgeCode

 ) ; 
 
 
// generating the bitmap 
 


	localparam logic [11:0] TRANSPARENT_ENCODING = 12'h000 ;// RGB value in the bitmap representing a transparent pixel  
	logic[0:31][0:63] object_colors = {
	64'b0000000000000000111111000011110011100011111100001110000000000000,
	64'b0000000000000001111111110011110011100011111110001110000000000000,
	64'b0000000000000001110011110011110011100011111110001110000000000000,
	64'b0000000000000001110011110011110011100011101110001110000000000000,
	64'b0000000000000001111000000011110111100011101110001110000000000000,
	64'b0000000000000001111111100011111111100011101111001110000000000000,
	64'b0000000000000000011111110011111111100111101111001110000000000000,
	64'b0000000000000000000011110011110011100111111111001110000000000000,
	64'b0000000000000001110011110011110011100111111111001110000000000000,
	64'b0000000000000001111011110011110011100111000111001110000000000000,
	64'b0000000000000000111111100011110011101111000111001110000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0011111100011110011111110000111110000111100000111111101111111100,
	64'b0011111110011110011111110011111111100111100000111111101111111110,
	64'b0000011111011110011110000011110111100111100000111100001111001111,
	64'b0000011111011110011110000011110111100111100000111000001111001111,
	64'b0000111110011110011110000011110000000111100000111100001111001111,
	64'b0001111100011110011111110011110000000111100000111111001111111110,
	64'b0001111000011110011111110011110111100111100000111111001111111110,
	64'b0011110000011110011110000011110111100111100000111000001111001111,
	64'b0111110000011110011110000011110111100111100000111000001111001111,
	64'b1111100000011110011110000011110111100111100000111100001111001111,
	64'b0111111110011110011111111011111111100111111110111111101111001111,
	64'b0011111110011110011111111000111110000111111110111111101111001111};	 
	//////////--------------------------------------------------------------------------------------------------------------= 
	//hit bit map has one bit per edge:  hit_colors[3:0] =   {Left, Top, Right, Bottom}	 
	//there is one bit per edge, in the corner two bits are set  
	 logic [0:3] [0:3] [3:0] hit_colors = 
				{16'h746,     
				16'h762,    
				16'h72, 
				16'h73}; 
	 // pipeline (ff) to get the pixel color from the array 	 
	//////////--------------------------------------------------------------------------------------------------------------= 
	always_ff@(posedge clk or negedge resetN) 
	begin 
		if(!resetN) begin 
			RGBout <=	3'h7; 
			HitEdgeCode <= 4'h0; 
		end 
		else begin 
			RGBout <= TRANSPARENT_ENCODING ; // default  
			HitEdgeCode <= 4'h0; 
	 
			if (InsideRectangle == 1'b1 ) 
			begin // inside an external bracket  
				HitEdgeCode <= hit_colors[offsetY >> 6][offsetX >> 6 ]; // get hitting edge from the colors table
				RGBout <= object_colors[offsetY][offsetX]? 12'hFFF : 12'h000 ;
			end
			else begin
				RGBout <= TRANSPARENT_ENCODING ; // default  
			end 		
			 
		end 
	end 
	 
	//////////--------------------------------------------------------------------------------------------------------------= 
	// decide if to draw the pixel or not 
	assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   




endmodule 
