module background(
	input	logic	clk,
	input	logic	resetN,
	input 	[10:0] 	pixelX,
	input 	[10:0]	pixelY,
	output 	[11:0] 	background_RGB
	
	
);



logic[0:31][0:31][1:0] object_colors = {
{2'h3,2'h3,2'h3,2'h3,2'h1,2'h2,2'h2,2'h3,2'h3,2'h3,2'h1,2'h3,2'h3,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h3,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h3,2'h3,2'h3,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h3,2'h3,2'h3,2'h1,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h3,2'h3,2'h3,2'h1,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h3,2'h3,2'h3,2'h2,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h3,2'h3,2'h2,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h3,2'h3,2'h2,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h3,2'h2,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h2,2'h2,2'h1},
{2'h3,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h1,2'h1,2'h2,2'h2,2'h2},
{2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h1,2'h2,2'h2,2'h3},
{2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h1,2'h2,2'h2,2'h2},
{2'h1,2'h1,2'h2,2'h2,2'h2,2'h2,2'h2,2'h1,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h2,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1},
{2'h3,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1},
{2'h3,2'h3,2'h3,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1},
{2'h3,2'h3,2'h3,2'h3,2'h1,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1},
{2'h3,2'h3,2'h3,2'h3,2'h3,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1},
{2'h3,2'h3,2'h3,2'h3,2'h3,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1},
{2'h3,2'h3,2'h3,2'h3,2'h1,2'h1,2'h1,2'h1,2'h2,2'h2,2'h2,2'h2,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1},
{2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h3,2'h2,2'h2,2'h2,2'h2,2'h3,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2},
{2'h2,2'h2,2'h3,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2},
{2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h1,2'h1,2'h1,2'h2,2'h2,2'h1,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h1,2'h1,2'h1,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2,2'h2},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h3,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h2,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h3,2'h3,2'h3,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h1,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h3,2'h3,2'h3,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h1,2'h2,2'h1},
{2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h1,2'h3,2'h1,2'h1,2'h1}};	
	
always_ff@(posedge clk or negedge resetN)
	begin
		if(!resetN) begin
			background_RGB <=	12'h000;

		end
		else begin
			case (object_colors[pixelY[7:0]][pixelX[7:0]])
				2'h1: background_RGB <= 12'hc60;
				2'h2: background_RGB <= 12'hFFC;
				2'h3: background_RGB <= 12'h630;
			endcase
		end
				
	end
	
endmodule
