
 module win_screen_bitmap (

	input	logic	clk, 
	input	logic	resetN, 
	input logic	[10:0] offsetX,// offset from top left  position 
	input logic	[10:0] offsetY, 
	input	logic	InsideRectangle, //input that the pixel is within a bracket 

	output	logic	drawingRequest, //output that the pixel should be dispalyed 
	output	logic	[11:0] RGBout,  //rgb value from the bitmap 
	output	logic	[3:0] HitEdgeCode

 ) ; 
 
 
// generating the bitmap 
 


	localparam logic [11:0] TRANSPARENT_ENCODING = 12'h000 ;// RGB value in the bitmap representing a transparent pixel  
	logic[0:255][0:255] object_colors = {
		256'b0011111111111111111111111111111111000000000000000000111111111111111111111111111110000000000000000001111111111111111111111111111111111110000000000000000000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0011111111111111111111111111111111000000000000000001111111111111111111111111111110000000000000000011111111111111111111111111111111111111000000000000000000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0011111111111111111111111111111111000000000000000011111111111111111111111111111110000000000000000111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0001111111111111111111111111111111000000000000000011111111111111111111111111111100000000000001111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000111111111111111111111111111111000000000000000011111111111111111111111111111000000000000001111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000111111111111111111111111111111000000000000000011111111111111111111111111111000000000000111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000111111111111111111111111111111000000000000000011111111111111111111111111111000000000011111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000111111111111111111111111111111100000000000000111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000011111111111111111111111111111110000000000001111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000001111111111111111111111111111110000000000001111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000001111111111111111111111111111110000000000001111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000111111111111111111111111111110000000000001111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000011111111111111111111111111110000000000001111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000011111111111111111111111111111000000000001111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000011111111111111111111111111111100000000011111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000001111111111111111111111111111100000000111111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000111111111111111111111111111100000000111111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000111111111111111111111111111100000000111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000111111111111111111111111111100000000111111111111111111111111111000000001111111111111111111111111111111000000001111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000111111111111111111111111111110000000111111111111111111111111111000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000011111111111111111111111111111000001111111111111111111111111111000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000001111111111111111111111111111000011111111111111111111111111110000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000001111111111111111111111111111000011111111111111111111111111100000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000001111111111111111111111111111000011111111111111111111111111100000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000111111111111111111111111111000011111111111111111111111111000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000011111111111111111111111111000011111111111111111111111110000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000011111111111111111111111111100111111111111111111111111110000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000011111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000011111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000001111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000011111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000001111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000001111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000001111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000001111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000011111111111111111111111111111111111111111111000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000011111111111111111111111111111111111111111111000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000011111111111111111111111111111111111111111111000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000001111111111111111111111111111111111111111110000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000111111111111111111111111111111111111111100000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000111111111111111111111111111111111111111100000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000111111111111111111111111111111111111111100000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000111111111111111111111111111111111111111100000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000011111111111111111111111111111111111111000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000001111111111111111111111111111111111110000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000001111111111111111111111111111111111110000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000001111111111111111111111111111111111110000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000111111111111111111111111111111111100000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111111000000001111111111111111111111111111111110000000000001111111111111111111111111111110000000011111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111100000000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000000001111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000000001111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000000000011111111111111111111111111111111111111111111111111111100000000000000000000000000000011111111111111111111111111111111111111111111111111111000000000000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111111111111111111000000000000000000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111111111111111111000000000000000000000000000000000000,
		256'b0000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		256'b1111111111111111111111111111110000000000000011111111111111000000000000011111111111111111111111111110000000000000000000011111111111111111111111111111111111111000000000000000000000000000011111111111111111111111111100000000000000001111111111111111111111111111,
		256'b1111111111111111111111111111110000000000000011111111111111000000000000011111111111111111111111111110000000000000000001111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111100000000000000001111111111111111111111111111,
		256'b1111111111111111111111111111110000000000000011111111111111000000000000011111111111111111111111111110000000000000000001111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111100000000000000001111111111111111111111111111,
		256'b0111111111111111111111111111110000000000000011111111111111000000000000111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111100000000000000001111111111111111111111111111,
		256'b0011111111111111111111111111110000000000000011111111111111000000000001111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111100000000000000001111111111111111111111111111,
		256'b0011111111111111111111111111110000000000000111111111111111000000000001111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111110000000000000001111111111111111111111111111,
		256'b0011111111111111111111111111111000000000001111111111111111000000000001111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111000000000000001111111111111111111111111111,
		256'b0011111111111111111111111111111100000000001111111111111111000000000001111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111000000000000001111111111111111111111111111,
		256'b0011111111111111111111111111111100000000001111111111111111100000000001111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111000000000000001111111111111111111111111111,
		256'b0011111111111111111111111111111100000000001111111111111111110000000001111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111100000000000001111111111111111111111111111,
		256'b0001111111111111111111111111111100000000001111111111111111110000000001111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111110000000000001111111111111111111111111111,
		256'b0000111111111111111111111111111100000000001111111111111111110000000001111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111110000000000001111111111111111111111111111,
		256'b0000111111111111111111111111111100000000001111111111111111110000000001111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111110000000000001111111111111111111111111111,
		256'b0000111111111111111111111111111100000000001111111111111111110000000001111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111110000000000001111111111111111111111111111,
		256'b0000111111111111111111111111111100000000001111111111111111110000000011111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111000000000001111111111111111111111111111,
		256'b0000111111111111111111111111111100000000001111111111111111110000000111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111100000000001111111111111111111111111111,
		256'b0000111111111111111111111111111100000000001111111111111111110000000111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111100000000001111111111111111111111111111,
		256'b0000111111111111111111111111111110000000011111111111111111110000000111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111100000000001111111111111111111111111111,
		256'b0000111111111111111111111111111111000000111111111111111111110000000111111111111111111111111111110000000111111111111111111111111111111100000000111111111111111111111111111111100000000000011111111111111111111111111111111110000000001111111111111111111111111111,
		256'b0000011111111111111111111111111111000000111111111111111111110000000111111111111111111111111111100000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111000000001111111111111111111111111111,
		256'b0000001111111111111111111111111111000000111111111111111111111000000111111111111111111111111111100000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111000000001111111111111111111111111111,
		256'b0000001111111111111111111111111111000000111111111111111111111100000111111111111111111111111111100000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111000000001111111111111111111111111111,
		256'b0000001111111111111111111111111111000000111111111111111111111100000111111111111111111111111111100000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111000000001111111111111111111111111111,
		256'b0000001111111111111111111111111111000000111111111111111111111100000111111111111111111111111111100000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111000000001111111111111111111111111111,
		256'b0000001111111111111111111111111111000000111111111111111111111100001111111111111111111111111111100000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111100000001111111111111111111111111111,
		256'b0000001111111111111111111111111111000000111111111111111111111100011111111111111111111111111111100000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111110000001111111111111111111111111111,
		256'b0000001111111111111111111111111111000000111111111111111111111100011111111111111111111111111111100000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111110000001111111111111111111111111111,
		256'b0000001111111111111111111111111111100000111111111111111111111100011111111111111111111111111111000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111110000001111111111111111111111111111,
		256'b0000000111111111111111111111111111110000111111111111111111111100011111111111111111111111111110000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111110000001111111111111111111111111111,
		256'b0000000011111111111111111111111111110000111111111111111111111100011111111111111111111111111110000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111000001111111111111111111111111111,
		256'b0000000011111111111111111111111111110001111111111111111111111100011111111111111111111111111110000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111100001111111111111111111111111111,
		256'b0000000011111111111111111111111111110011111111111111111111111100011111111111111111111111111110000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111100001111111111111111111111111111,
		256'b0000000011111111111111111111111111110011111111111111111111111100011111111111111111111111111110000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111100001111111111111111111111111111,
		256'b0000000011111111111111111111111111110011111111111111111111111110011111111111111111111111111110000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111110001111111111111111111111111111,
		256'b0000000011111111111111111111111111110011111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111001111111111111111111111111111,
		256'b0000000011111111111111111111111111110011111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111001111111111111111111111111111,
		256'b0000000011111111111111111111111111110011111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111001111111111111111111111111111,
		256'b0000000001111111111111111111111111110011111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111001111111111111111111111111111,
		256'b0000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000011111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000001111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000001111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000001111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000001111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000001111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000001111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000001111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000001111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000000111111111111111111111111111111111111100111111111111111111111111111111111110000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111,
		256'b0000000000000011111111111111111111111111111111111100111111111111111111111111111111111110000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111001111111111111111111111111111111111111111,
		256'b0000000000000011111111111111111111111111111111111100111111111111111111111111111111111110000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111001111111111111111111111111111111111111111,
		256'b0000000000000011111111111111111111111111111111111100111111111111111111111111111111111110000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111001111111111111111111111111111111111111111,
		256'b0000000000000011111111111111111111111111111111111100111111111111111111111111111111111110000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111001111111111111111111111111111111111111111,
		256'b0000000000000011111111111111111111111111111111111100111111111111111111111111111111111110000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000111111111111111111111111111111111111111,
		256'b0000000000000011111111111111111111111111111111111100111111111111111111111111111111111100000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000011111111111111111111111111111111111111,
		256'b0000000000000011111111111111111111111111111111111100111111111111111111111111111111111000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000011111111111111111111111111111111111111,
		256'b0000000000000011111111111111111111111111111111111000111111111111111111111111111111111000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000011111111111111111111111111111111111111,
		256'b0000000000000001111111111111111111111111111111110000111111111111111111111111111111111000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000011111111111111111111111111111111111111,
		256'b0000000000000000111111111111111111111111111111110000111111111111111111111111111111111000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000011111111111111111111111111111111111111,
		256'b0000000000000000111111111111111111111111111111110000011111111111111111111111111111111000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000001111111111111111111111111111111111111,
		256'b0000000000000000111111111111111111111111111111110000001111111111111111111111111111111000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000000111111111111111111111111111111111111,
		256'b0000000000000000111111111111111111111111111111110000001111111111111111111111111111111000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000000111111111111111111111111111111111111,
		256'b0000000000000000111111111111111111111111111111110000001111111111111111111111111111111000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000000111111111111111111111111111111111111,
		256'b0000000000000000111111111111111111111111111111110000001111111111111111111111111111110000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000000011111111111111111111111111111111111,
		256'b0000000000000000111111111111111111111111111111110000001111111111111111111111111111100000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000000001111111111111111111111111111111111,
		256'b0000000000000000111111111111111111111111111111110000001111111111111111111111111111100000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000000001111111111111111111111111111111111,
		256'b0000000000000000011111111111111111111111111111110000001111111111111111111111111111100000000000000000000111111111111111111111111111111000000000011111111111111111111111111111100000000000011111111111111111111111111111000000001111111111111111111111111111111111,
		256'b0000000000000000001111111111111111111111111111110000001111111111111111111111111111100000000000000000000111111111111111111111111111111100000000111111111111111111111111111111100000000000011111111111111111111111111111000000001111111111111111111111111111111111,
		256'b0000000000000000001111111111111111111111111111110000001111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111000000000111111111111111111111111111111111,
		256'b0000000000000000001111111111111111111111111111100000001111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111000000000011111111111111111111111111111111,
		256'b0000000000000000001111111111111111111111111111000000001111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111000000000011111111111111111111111111111111,
		256'b0000000000000000001111111111111111111111111111000000001111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111000000000011111111111111111111111111111111,
		256'b0000000000000000001111111111111111111111111111000000000111111111111111111111111111000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111000000000001111111111111111111111111111111,
		256'b0000000000000000001111111111111111111111111111000000000011111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111000000000000111111111111111111111111111111,
		256'b0000000000000000000111111111111111111111111111000000000011111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111000000000000111111111111111111111111111111,
		256'b0000000000000000000011111111111111111111111111000000000011111111111111111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111000000000000111111111111111111111111111111,
		256'b0000000000000000000011111111111111111111111111000000000011111111111111111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111000000000000111111111111111111111111111111,
		256'b0000000000000000000011111111111111111111111111000000000011111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111000000000000111111111111111111111111111111,
		256'b0000000000000000000011111111111111111111111111000000000011111111111111111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111000000000000011111111111111111111111111111,
		256'b0000000000000000000011111111111111111111111111000000000011111111111111111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111000000000000001111111111111111111111111111,
		256'b0000000000000000000011111111111111111111111111000000000011111111111111111111111110000000000000000000000000000000011111111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111000000000000001111111111111111111111111111,
		256'b0000000000000000000011111111111111111111111110000000000011111111111111111111111100000000000000000000000000000000000111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111000000000000001111111111111111111111111111,
		256'b0000000000000000000011111111111111111111111100000000000011111111111111111111111000000000000000000000000000000000000111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111000000000000001111111111111111111111111111,
		256'b0000000000000000000001111111111111111111111100000000000011111111111111111111111000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111000000000000000111111111111111111111111111,
		256'b0000000000000000000000111111111111111111111100000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000011111111111111111111111111111000000000000000011111111111111111111111111,
		256'b0000000000000000000000111111111111111111111100000000000000111111111111111111111000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000011111111111111111111111111111000000000000000011111111111111111111111111};
	 
	//////////--------------------------------------------------------------------------------------------------------------= 
	//hit bit map has one bit per edge:  hit_colors[3:0] =   {Left, Top, Right, Bottom}	 
	//there is one bit per edge, in the corner two bits are set  
	 logic [0:3] [0:3] [3:0] hit_colors = 
				{16'h746,     
				16'h762,    
				16'h72, 
				16'h73}; 
	 // pipeline (ff) to get the pixel color from the array 	 
	//////////--------------------------------------------------------------------------------------------------------------= 
	always_ff@(posedge clk or negedge resetN) 
	begin 
		if(!resetN) begin 
			RGBout <=	3'h7; 
			HitEdgeCode <= 4'h0; 
		end 
		else begin 
			RGBout <= TRANSPARENT_ENCODING ; // default  
			HitEdgeCode <= 4'h0; 
	 
			if (InsideRectangle == 1'b1 ) 
			begin // inside an external bracket  
				HitEdgeCode <= hit_colors[offsetY >> 6][offsetX >> 6 ]; // get hitting edge from the colors table
				RGBout <= object_colors[offsetY][offsetX]? 12'hFFF : 12'h000 ;
			end
			else begin
				RGBout <= TRANSPARENT_ENCODING ; // default  
			end 		
			 
		end 
	end 
	 
	//////////--------------------------------------------------------------------------------------------------------------= 
	// decide if to draw the pixel or not 
	assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   




endmodule 
