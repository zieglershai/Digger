
module	player_life_bitmap	(	
	input	logic	clk,
	input	logic	resetN,
	input logic	[10:0] offsetX,// offset from top left  position 
	input logic	[10:0] offsetY,
	input	logic	InsideRectangle, //input that the pixel is within a bracket 
	input logic playGame,
	input logic player_died,

	output	logic	drawingRequest, //output that the pixel should be dispalyed 
	output	logic	[11:0] RGBout,  //rgb value from the bitmap 
	output	logic no_lives

 ) ;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 5;  // 2^4 = 16
localparam  int OBJECT_NUMBER_OF_X_BITS = 5;  // 2^6 = 64


localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_HEIGHT_Y_DIVIDER = OBJECT_NUMBER_OF_Y_BITS - 2; //how many pixel bits are in every collision pixel
localparam  int OBJECT_WIDTH_X_DIVIDER =  OBJECT_NUMBER_OF_X_BITS - 2;

// generating a smiley bitmap

localparam logic [11:0] TRANSPARENT_ENCODING = 12'h000 ;// RGB value in the bitmap representing a transparent pixel 


logic unsigned [0:2] initial_life = { 1'b1, 1'b1, 1'b1}; //fukcer
logic unsigned [0:2] MazeBiMapMask;



logic [0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1][11:0] object_colors = {
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf90,12'hf90,12'hf90,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'hf90,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'hf90,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'hf00,12'hf00,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'hf00,12'hf00,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000}
	 };

//////////--------------------------------------------------------------------------------------------------------------=
//hit bit map has one bit per edge:  hit_colors[3:0] =   {Left, Top, Right, Bottom}	
//there is one bit per edge, in the corner two bits are set  


 

// pipeline (ff) to get the pixel color from the array 	 

//////////--------------------------------------------------------------------------------------------------------------=
	always_ff@(posedge clk  or negedge resetN)
	begin
		if(!resetN) begin
			MazeBiMapMask <= initial_life;
			no_lives <= 0;

		end
		


		else begin
			 /// for each collosion delete one life
			if (player_died) begin
				if (MazeBiMapMask[2])
					MazeBiMapMask[2] <= 0;
				else if (MazeBiMapMask[1])
					MazeBiMapMask[1] <= 0;
				/*else if (MazeBiMapMask[0])
					MazeBiMapMask[0] <= 0;
				*/
				else
					no_lives <= 1;
			end
				
		end
			
	end

//////////--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
	assign drawingRequest = MazeBiMapMask[offsetX[8:5]] && object_colors[offsetY][offsetX] != TRANSPARENT_ENCODING;  // in the area and have enough life and ligtehn pixel
	assign RGBout = object_colors[offsetY][offsetX];

endmodule