module score_bit_map	(	
	input		logic	clk,
	input		logic	resetN,
	input		logic	startOfFrame,
	input 	logic	[10:0] offsetX,// offset from top left  position 
	input 	logic	[10:0] offsetY,
	input		logic	InsideRectangle, //input that the pixel is within a bracket 
	input 	logic	player_eat_gold, // points to add
	input 	logic player_eat_dimond,
	
	output	logic				drawingRequest, //output that the pixel should be dispalyed 
	output	logic	[11:0]		RGBout

);



wire logic[4:0]  hunderes, thousands;
bit [0:9] [0:31] [0:15] number_bitmap  = {


{
// 0

	16'b0000111111110000,
	16'b0001111111111000,
	16'b0011111111111100,
	16'b0111111111111110,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b0111111111111110,
	16'b0011111111111100,
	16'b0001111111111000,
	16'b0000111111110000},
			
// 00
			
{
	16'b0000111111111111,
	16'b0000111111111111,
	16'b0000111111111111,
	16'b0000111111111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111,
	16'b0000000011111111},
		
// 11
{
	16'b0000111111110000,
	16'b0001111111111000,
	16'b0011111111111100,
	16'b0111111111111110,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b0000000000111111,
	16'b0000000001111111,
	16'b0000000011111111,
	16'b0000000111111111,
	16'b0000001111111100,
	16'b0000001111111100,
	16'b0000011111111100,
	16'b0000111111111000,
	16'b0001111111110000,
	16'b0011111111100000,
	16'b0011111111000000,
	16'b0011111110000000,
	16'b0111111100000000,
	16'b1111110000000000,
	16'b1111110000000000,
	16'b1111110000000000,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111111111111111},
	
// 3
{	
	16'b0000111111110000,
	16'b0001111111111000,
	16'b0011111111111100,
	16'b0111111111111110,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b0000000000111111,
	16'b0000000001111111,
	16'b0000000011111110,
	16'b0000000111111100,
	16'b0000001111110000,
	16'b0000001111110000,
	16'b0000001111110000,
	16'b0000001111110000,
	16'b0000000000111100,
	16'b0000000000111100,
	16'b0000000000111111,
	16'b0000000000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b0111111111111110,
	16'b0011111111111100,
	16'b0001111111111000,
	16'b0000111111110000},
			
// 4
																			
{
	16'b0000000011110000,
	16'b0000000011110000,
	16'b0000000011110000,
	16'b0000000111110000,
	16'b0000001111110000,
	16'b0000001111110000,
	16'b0000001111110000,
	16'b0000011111110000,
	16'b0000111111110000,
	16'b0000111111110000,
	16'b0000111111110000,
	16'b0001111111110000,
	16'b0011110011110000,
	16'b0011110011110000,
	16'b0011110011110000,
	16'b0011110011110000,
	16'b0011000011110000,
	16'b0111000011110000,
	16'b1111000011110000,
	16'b1111000011110000,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b0111111111111110,
	16'b0011111111111100,
	16'b0000000111111000,
	16'b0000000011110000,
	16'b0000000011110000,
	16'b0000000011110000,
	16'b0000000011110000,
	16'b0000000011110000},
			
			
// 5
																			
{
	16'b1111111111111100,
	16'b1111111111111100,
	16'b1111111111111100,
	16'b1111111111111100,
	16'b1111111111111100,
	16'b1111111111111100,
	16'b1111110000000000,
	16'b1111110000000000,
	16'b1111110000000000,
	16'b1111110000000000,
	16'b1111110000000000,
	16'b1111110000000000,
	16'b1111111111110000,
	16'b1111111111111000,
	16'b0111111111111100,
	16'b0011111111111110,
	16'b0001111111111111,
	16'b0000111111111111,
	16'b0000000000111111,
	16'b0000000000111111,
	16'b0000000000111111,
	16'b0000000000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b0011111111111110,
	16'b0011111111111100,
	16'b0001111111111000,
	16'b0000111111110000},
			
			
// 6
																			
{
	16'b0000111111110000,
	16'b0000111111111000,
	16'b0011111111111100,
	16'b0011111111111110,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000000000,
	16'b1111110000000000,
	16'b1111110000000000,
	16'b1111110000000000,
	16'b1111111111111100,
	16'b1111111111111110,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b0111111111111110,
	16'b0011111111111100,
	16'b0001111111111000,
	16'b0000111111110000},
			
// 7
																			
{
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b0000000000111100,
	16'b0000000000111100,
	16'b0000000011111100,
	16'b0000000011111100,
	16'b0000000011111100,
	16'b0000000111111100,
	16'b0000001111111000,
	16'b0000001111110000,
	16'b0000001111110000,
	16'b0000001111110000,
	16'b0000001111110000,
	16'b0000011111110000,
	16'b0000111111100000,
	16'b0000111111000000,
	16'b0000111111000000,
	16'b0000111111000000,
	16'b0000111111000000,
	16'b0001111111000000,
	16'b0011111110000000,
	16'b0011111100000000,
	16'b0011111100000000,
	16'b0011111100000000,
	16'b0011111100000000,
	16'b0011111100000000
},
			
// 16
																			
{
	16'b0000111111110000,
	16'b0001111111111000,
	16'b0011111111111100,
	16'b0111111111111110,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b0111111111111110,
	16'b0011111111111100,
	16'b0011111111111000,
	16'b0011111111111000,
	16'b0011111111111100,
	16'b0111111111111100,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b0111111111111110,
	16'b0011111111111100,
	16'b0001111111111000,
	16'b0000111111110000},
			
// 9
																			
{
	16'b0000111111110000,
	16'b0001111111111000,
	16'b0011111111111100,
	16'b0111111111111110,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b0011111111111111,
	16'b0011111111111111,
	16'b0000000000111111,
	16'b0000000000111111,
	16'b0000000000111111,
	16'b0000000000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111110000111111,
	16'b1111111111111111,
	16'b1111111111111111,
	16'b0111111111111110,
	16'b0011111111111100,
	16'b0001111111111000,
	16'b0000111111110000}


};


	always_ff@(posedge clk or negedge resetN)
	begin
		if(!resetN) begin
			hunderes <= 5'b0;
			thousands <= 5'b0;
		end
		else begin
			if (player_eat_gold) begin
				if (hunderes == 5'd9) begin
					thousands <= thousands + 5'd1;
					hunderes  <= 5'b1;
				end
				else if (hunderes == 5'd8) begin
					thousands <= thousands + 5'd1;
					hunderes  <= 5'b0;
				end
				else begin
					hunderes  <= hunderes +  5'd2;
				end
			end
			if (player_eat_dimond)begin
				if (hunderes == 5'd9) begin
					thousands <= thousands + 5'd1;
					hunderes  <= 5'b0;
				end
				else begin
					hunderes  <= hunderes +  5'd1;
				end
			end
		end
	end

	always_comb begin
		if (offsetX[7:4] == 4'd0)begin
			RGBout = number_bitmap[thousands][offsetY[4:0]][offsetX[3:0]]? 12'h000 : 12'hFFF ; // this is a fixed color
		end
		else if (offsetX[7:4] == 4'd1)begin
			RGBout = number_bitmap[hunderes][offsetY[4:0]][offsetX[3:0]]? 12'h000 : 12'hFFF  ; // this is a fixed color
		end
		else begin
			RGBout = number_bitmap[5'd0][offsetY[4:0]][offsetX[3:0]]? 12'h000 : 12'hFFF  ; // this is a fixed color
		end
	end
	
	
	
	assign drawingRequest =  InsideRectangle & (!RGBout[0]); 

endmodule 