
module	alien_bitmap	(	
					input	logic	clk,
					input	logic	resetN,
					input startOfFrame,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input	logic	playerHit, //input that the pixel is within a bracket 

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[11:0] RGBout,  //rgb value from the bitmap 
					output	logic	[3:0] HitEdgeCode //one bit per edge 
 ) ;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 5;  // 2^4 = 16
localparam  int OBJECT_NUMBER_OF_X_BITS = 5;  // 2^6 = 64


localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_HEIGHT_Y_DIVIDER = OBJECT_NUMBER_OF_Y_BITS - 2; //how many pixel bits are in every collision pixel
localparam  int OBJECT_WIDTH_X_DIVIDER =  OBJECT_NUMBER_OF_X_BITS - 2;

// generating a smiley bitmap

localparam logic [11:0] TRANSPARENT_ENCODING = 12'hFFF ;// RGB value in the bitmap representing a transparent pixel 

logic [2:0][0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1][11:0] object_colors = {
{
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h000,12'h000,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h900,12'hFF3,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h900,12'h900,12'hFF3,12'h900,12'hBF6,12'h000,12'h000,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h900,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'h900,12'hFF3,12'h8F0,12'hFF3,12'h8F0,12'h8F0,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'hFF3,12'h8F0,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'h000,12'hFF3,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'h000,12'hFF3,12'hFF3,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'h900,12'h8F0,12'hFF3,12'hBF6,12'hBF6,12'h8F0,12'h8F0,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'h900,12'hFF3,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h900,12'h900,12'hFF3,12'h8F0,12'hFF3,12'hBF6,12'hBF6,12'hFF3,12'h8F0,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h900,12'hFF3,12'hFF3,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hBF6,12'hBF6,12'hBF6,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h900,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h900,12'hFF3,12'h8F0,12'h8F0,12'hFF3,12'hBF6,12'hBF6,12'hBF6,12'hBF6,12'h8F0,12'hFF3,12'hFF3,12'hFF3,12'h900,12'hFF3,12'hFF3,12'h900,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hFF3,12'h900,12'hFF3,12'hFF3,12'h8F0,12'hFF3,12'h8F0,12'hFF3,12'hFF3,12'h8F0,12'hBF6,12'hBF6,12'hBF6,12'hFF3,12'h8F0,12'hFF3,12'hFF3,12'h8F0,12'hFF3,12'hFF3,12'hBF6,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h000,12'h000,12'hFF3,12'h8F0,12'h8F0,12'hFF3,12'hBF6,12'hBF6,12'hBF6,12'h8F0,12'hBF6,12'h8F0,12'h8F0,12'hBF6,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hBF6,12'h000,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h000,12'h000,12'h000,12'hBF6,12'h8F0,12'hFF3,12'hBF6,12'hBF6,12'h8F0,12'h000,12'h000,12'hBF6,12'h8F0,12'hBF6,12'hBF6,12'h8F0,12'hBF6,12'h000,12'h000,12'h000,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h000,12'h000,12'h000,12'hBF6,12'hFF3,12'h8F0,12'hBF6,12'h8F0,12'h8F0,12'h000,12'h000,12'h000,12'hBF6,12'hBF6,12'hBF6,12'h8F0,12'hBF6,12'h000,12'h000,12'h000,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h000,12'h000,12'h000,12'hFF3,12'hBF6,12'h8F0,12'h8F0,12'h8F0,12'h000,12'h000,12'h000,12'h000,12'hBF6,12'hBF6,12'h8F0,12'hBF6,12'hBF6,12'hFF3,12'h000,12'h000,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h000,12'h900,12'h900,12'h900,12'hFF3,12'h8F0,12'h8F0,12'hFF3,12'h000,12'h000,12'h000,12'h000,12'h000,12'h8F0,12'hBF6,12'hBF6,12'h900,12'h900,12'h900,12'h000,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h900,12'hFF3,12'h900,12'h000,12'hFF3,12'hBF6,12'h8F0,12'h8F0,12'hBF6,12'h000,12'h000,12'h000,12'hBF6,12'hBF6,12'hBF6,12'h000,12'hFF3,12'hFC9,12'h900,12'h000,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h900,12'hFB0,12'h000,12'h000,12'h000,12'h000,12'hBF6,12'h8F0,12'hFF3,12'h000,12'h000,12'h000,12'hBF6,12'hBF6,12'h000,12'h000,12'hFF3,12'hFF3,12'hFC9,12'h000,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'h900,12'h900,12'h000,12'h000,12'h000,12'h000,12'hBF6,12'h8F0,12'hFF3,12'hBF6,12'h000,12'hBF6,12'hBF6,12'hBF6,12'h000,12'h000,12'h000,12'h900,12'hFC9,12'h900,12'h900,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'h900,12'hFC9,12'hF80,12'h900,12'h000,12'h000,12'h000,12'h000,12'h8F0,12'h8F0,12'h8F0,12'hBF6,12'hBF6,12'hBF6,12'h000,12'h000,12'h000,12'h000,12'h000,12'hFC9,12'h900,12'h900,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFC9,12'hFB0,12'hF80,12'h900,12'h000,12'h000,12'h000,12'h000,12'h000,12'h8F0,12'hBF6,12'h8F0,12'hBF6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hFB0,12'hFB0,12'h900,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'h000,12'h900,12'hFC9,12'hFB0,12'hF80,12'hF80,12'hF80,12'h900,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hFC9,12'hF80,12'h900,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'h900,12'hFF3,12'hFC9,12'hFC9,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hFB0,12'hFB0,12'hF80,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'h900,12'hFF3,12'hFC9,12'hFC9,12'hFB0,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h900,12'hFC9,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'h900,12'hFC9,12'hFC9,12'hFB0,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'h900,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hFC9,12'hFB0,12'hFB0,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hFC9,12'hFB0,12'hFC9,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hFC9,12'hFB0,12'hFC9,12'hFB0,12'hF80,12'hF80,12'hF80,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h900,12'h900,12'hFC9,12'hFB0,12'hFB0,12'hF80,12'hF80,12'hF80,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h900,12'h900,12'h900,12'hFC9,12'h900,12'h900,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF}
	},
	
	{{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hFFC,12'hFF3,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFFF,12'hFF3,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'h900,12'h8F0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'h900,12'hFFF,12'h8F0,12'hFFF,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFFC,12'hFFC,12'hFFC,12'h900,12'hFFC,12'hFFC,12'hFFC,12'hFF3,12'hBF6,12'h8F0,12'hBF6,12'hBF6,12'hFFC,12'hFFC,12'hFFC,12'hF80,12'hFFC,12'hFFC,12'hFFC,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFC,12'hFFC,12'hFFC,12'h000,12'h000,12'h900,12'hFFC,12'hFFC,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'hBF6,12'hFFC,12'hFFC,12'h000,12'h000,12'hFFC,12'hFFC,12'hFFC,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFFC,12'hFFC,12'h000,12'h000,12'h900,12'hFFC,12'hFF3,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'hBF6,12'hBF6,12'hFFC,12'h000,12'h000,12'h900,12'hFFC,12'hFFC,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFC,12'hFFC,12'hFFC,12'hFFC,12'h900,12'hFFC,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'h900,12'h8F0,12'h000,12'hFFC,12'hFFC,12'hFFC,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFC,12'hFFC,12'h900,12'hFF3,12'hFF3,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hFF3,12'h900,12'hFFC,12'hFF3,12'hFFC,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h900,12'hBF6,12'hBF6,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hFF3,12'h900,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hBF6,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h000,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFFC,12'hFFC,12'hF80,12'h000,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFC,12'hFFC,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFC,12'hF80,12'hF80,12'h900,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFC,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hF80,12'hF80,12'h900,12'h900,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'h000,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'h900,12'hF80,12'hF80,12'hF80,12'h900,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'hFFF,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hF80,12'hFFC,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hFFC,12'hFFC,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'h900,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFC,12'hF80,12'hFFC,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h000,12'h000,12'h900,12'h900,12'h900,12'h900,12'h900,12'h900,12'h900,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFFC,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFC,12'hF80,12'hFFC,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'hF80,12'h900,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF}
	},
	{
	{12'hFFF,12'hFF3,12'h900,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hBF6,12'hFF3,12'hBF6,12'hBF6,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'h900,12'hBF6,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'h900,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hBF6,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hBF6,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h900,12'h000,12'h000,12'h000,12'hFF3,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'h000,12'hFF3,12'hFF3,12'hBF6,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h900,12'h000,12'h000,12'h000,12'hFF3,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'h000,12'hFF3,12'hFF3,12'hBF6,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h900,12'h000,12'h000,12'h000,12'hFF3,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'h000,12'h000,12'h000,12'hFF3,12'hBF6,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hBF6,12'hFF3,12'hFF3,12'h900,12'h000,12'h000,12'h000,12'hFF3,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hBF6,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hBF6,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hBF6,12'hBF6,12'hBF6,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hBF6,12'hBF6,12'hBF6,12'hBF6,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFF3,12'hFF3,12'hFF3,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFF3,12'hFF3,12'hFF3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h000,12'h000,12'h000,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h000,12'h000,12'h000,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFC9,12'h900,12'h900,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h000,12'h000,12'h000,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h900,12'h900,12'h900,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h000,12'h000,12'h000,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'h900,12'hFC9,12'hFC9,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'h900,12'hFC9,12'hFC9,12'h900,12'h900,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'h900,12'hFC9,12'hFB6,12'hFC9,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFC9,12'hFB6,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'hFFF,12'hFC9,12'hFB6,12'hFB6,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFC9,12'hFB6,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFC9,12'hFB6,12'hFB6,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFC9,12'hFC9,12'hFB6,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFC9,12'hFB6,12'hFB6,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFC9,12'hFB6,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8F0,12'h8F0,12'h8F0,12'h8F0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFC9,12'hFB6,12'hFB6,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFC9,12'hFB6,12'hFB6,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFC9,12'hFB6,12'hFB6,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFC9,12'hFB6,12'hFB6,12'hFC9,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFC9,12'hFB6,12'hFB6,12'hFC9,12'h900,12'h900,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'h900,12'hFC9,12'hFB6,12'hFB6,12'hFB6,12'hFB6,12'hFC9,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFC9,12'hFC9,12'hFB6,12'hFB6,12'hFC9,12'hFC9,12'hFC9,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFC9,12'hFB6,12'hFB6,12'hFB6,12'hFB6,12'hFB6,12'hFB6,12'hFC9,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFC9,12'hFB6,12'hFB6,12'hFB6,12'hFB6,12'hFB6,12'hFB6,12'hFC9,12'hFFF,12'hFFF,12'hFFF},
	{12'h900,12'hFC9,12'hFC9,12'hFC9,12'hFB6,12'hFB6,12'hFB6,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFC9,12'hFC9,12'hFC9,12'hFB6,12'hFB6,12'hFB6,12'hFB6,12'hFC9,12'hFC9,12'hFC9,12'h900,12'hFFF},
	{12'h900,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'h900,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h900,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'hFC9,12'h900,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
	{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF}
	}
	};

//////////--------------------------------------------------------------------------------------------------------------=
//hit bit map has one bit per edge:  hit_colors[3:0] =   {Left, Top, Right, Bottom}	
//there is one bit per edge, in the corner two bits are set  


logic [0:3] [0:3] [3:0] hit_colors = 
		  {16'hC446,     
			16'h8C62,    
			16'h8932,
			16'h9113};

 

// pipeline (ff) to get the pixel color from the array 	 


wire [8:0] counter;


//////////--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	12'h000;
		HitEdgeCode <= 4'h0;
		counter <= 9'b0;

	end
	else begin
		
		if (startOfFrame)begin
			counter <= counter + 9'b1;
		end
		if (InsideRectangle == 1'b1 ) begin
		 // inside an external bracket 
			HitEdgeCode <= hit_colors[offsetY >> OBJECT_HEIGHT_Y_DIVIDER][offsetX >> OBJECT_WIDTH_X_DIVIDER];	//get hitting edge from the colors table  
			if (counter[6:5] == 2'd3) begin
				RGBout <= object_colors[1][offsetY][offsetX];
			end
			else begin
				RGBout <= object_colors[counter[6:5]][offsetY][offsetX];
			end
		end  	
	end
		
end

//////////--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING && InsideRectangle) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   

endmodule