
module	player_bit_map	(	
					input	logic	clk,
					input	logic	resetN,
					input startOfFrame,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input	logic	playerHit, //input that the pixel is within a bracket 
					input	logic	[1:0] player_direction,
					input	logic	[2:0] image,			
					input logic player_awake,
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[11:0] RGBout,  //rgb value from the bitmap 
					output	logic	[3:0] HitEdgeCode //one bit per edge 
 ) ;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 5;  // 2^4 = 16
localparam  int OBJECT_NUMBER_OF_X_BITS = 5;  // 2^6 = 64


localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_HEIGHT_Y_DIVIDER = OBJECT_NUMBER_OF_Y_BITS - 2; //how many pixel bits are in every collision pixel
localparam  int OBJECT_WIDTH_X_DIVIDER =  OBJECT_NUMBER_OF_X_BITS - 2;

// generating a smiley bitmap

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel 

logic [0:1][0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [11:0] object_colors = {
	{{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf90,12'hf90,12'hf90,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'hf90,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'hf90,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'hf00,12'hf00,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'hf00,12'hf00,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000}},
	
	{{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'hf00,12'hf00,12'hf00,12'hf90,12'hf90,12'hf90,12'hf00,12'hf00,12'h0f6,12'hf00,12'hf00,12'h000,12'hf90,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'hf90,12'hf00,12'h0f6,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'hf90,12'hf00,12'h0f6,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'hf00,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h0f6,12'hf00,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000},
    {12'h000,12'hf00,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h0f6,12'hf00,12'hf00,12'hf00,12'hf00,12'h000,12'h000,12'h000,12'h000,12'hf00,12'hf00,12'hf00,12'h0f6,12'h0f6,12'h0f6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf00,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'hf00,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf00,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'hf00,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hf90,12'hf90,12'hf90,12'hf90,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
    {12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000}},
	 };
logic [0:3][0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [11:0] rip_colors = {

	 
	 {{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000}},

	 
	{{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'h4C6,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000}},

	{{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'hc94,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000},
	{12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94}},
	
	{{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'h000,12'h000,12'h4C6,12'h4C6,12'h4C6,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h4C6,12'h4C6,12'h000,12'h000},
	{12'hc94,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000},
	{12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'h000},
	{12'h000,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'h000,12'h000,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'hc94,12'h000,12'hc94,12'hc94,12'hc94}}
	
	
	 };
//////////--------------------------------------------------------------------------------------------------------------=
//hit bit map has one bit per edge:  hit_colors[3:0] =   {Left, Top, Right, Bottom}	
//there is one bit per edge, in the corner two bits are set  


logic [0:3] [0:3] [3:0] hit_colors = 
		  {16'hC446,     
			16'h8C62,    
			16'h8932,
			16'h9113};

 

// pipeline (ff) to get the pixel color from the array 	 


wire [7:0] counter;

//////////--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	12'h00;
		HitEdgeCode <= 4'h0;
		counter <= 8'h0;

	end
	else begin
		if (startOfFrame) begin
			counter <= counter + 8'h1;
		end
		else begin
			counter <= counter;
		end
		if (InsideRectangle == 1'b1 ) begin
		 // inside an external bracket 
			HitEdgeCode <= hit_colors[offsetY >> OBJECT_HEIGHT_Y_DIVIDER][offsetX >> OBJECT_WIDTH_X_DIVIDER];	//get hitting edge from the colors table  
			if (player_awake == 1'b1)begin
				if (player_direction == 2'b00) begin
					RGBout <= object_colors[counter[4]][offsetX][11'd32 - offsetY];
				end
				else if (player_direction == 2'b01) begin
					RGBout <= object_colors[counter[4]][offsetY][offsetX];

				end	
				else if (player_direction == 2'b10) begin
					RGBout <= object_colors[counter[4]][11'd32 - offsetX][offsetY];
				end
				else  begin
					RGBout <= object_colors[counter[4]][offsetY][11'd32 - offsetX];
				end	
			end
			else begin
				RGBout <= rip_colors [image][offsetY][offsetX];
			end
		end
		else begin
			RGBout <= TRANSPARENT_ENCODING;
		end

	end
		
end

//////////--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   

endmodule